**.subckt dc_res_temp
Vres Vcc GND 1.5
Vsil Vcc net1 0
Vppd Vcc net2 0
Vrh Vcc net3 0
XR1 GND net1 rsil w=0.5e-6 l=1.5e-6 m=1 b=0
XR2 GND net2 rppd w=0.5e-6 l=0.5e-6 m=1 b=0
XR3 GND net3 rhigh w=0.5e-6 l=0.5e-6 m=1 b=0
**** begin user architecture code

.include /foss/pdks/sg13g2/libs.tech/xyce/models/resistors.lib

.dc Vres 0 1.5 0.01
.PRINT  dc format=raw file=dc_res_temp.raw  I(Vsil) I(Vppd)  I(Vrh)

**** end user architecture code
**.ends
.GLOBAL GND
.end
