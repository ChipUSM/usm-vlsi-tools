** sch_path: TOP_ldo_cl_psrr.sch
**.subckt TOP_ldo_cl_psrr
V1 vcm_ldo1 vss 0.9
V5 vss GND 0
I0 vss iref_ldo1 5u
Cc net1 vss 10u m=1
Resr vout_ldo1 net1 2 m=1
Resr1 vout_ldo1 vss 12 m=1
Cc1 vout_ldo1 vss 50p m=1
Vs vdd_ldo1 vss 1.8 AC 1
x1 net2 net3 net4 net5 net6 net7 net8 vout_ldo1 net9 vdd_ldo1 net10 vcm_ldo1 net11 net12 iref_ldo1 net13 net14 net15 net16 net17  net18 vss net19 net20 net21 net22 net23 net24 TOP
**** begin user architecture code

.lib /opt/pdks/sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.lib /opt/pdks/sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ
.lib /opt/pdks/sg13g2/libs.tech/ngspice/models/cornerCAP.lib cap_typ

.option TEMP=27
.option warn=1

.control

pre_osdi /opt/pdks/sg13g2/libs.tech/ngspice/openvaf/psp103_nqs.osdi

** PSRR is defined as the change in input offset vs. change in power supply.
ac dec 100 1 10G
meas ac psrr find vdb(vout_ldo1) at=1

wrdata ngspice/psrr_1.data psrr
.endc

.GLOBAL GND


** sch_path: /home/ac3e/Documents/ihp_design/xschem/top/TOP.sch
.subckt TOP 28 22 23 24 26 27 25 1 21 2 20 3 19 18 4 5 17 6 16 15 7 8 9 10 11 12 13 14
*.PININFO 1:B 2:B 3:B 4:B 5:B 6:B 7:B 21:B 20:B 19:B 18:B 17:B 16:B 15:B 14:B 13:B 12:B 11:B 10:B 9:B 8:B 22:B 23:B 24:B 25:B 26:B
*+ 27:B 28:B
x1 2 1 4 3 8 ldo_closeloop
x2 28 25 26 27 8 24 23 ldo_openloop
x3 19 22 20 pass_transistor
x4 18 16 15 14 8 17 ota
.ends

* expanding   symbol:  xschem/ldo/ldo_closeloop.sym # of pins=5
** sym_path: /home/ac3e/Documents/ihp_design/xschem/ldo/ldo_closeloop.sym
** sch_path: /home/ac3e/Documents/ihp_design/xschem/ldo/ldo_closeloop.sch
.subckt ldo_closeloop ldo_in ldo_out iref vref vss
*.PININFO vss:B ldo_in:B ldo_out:O iref:I vref:I
XM1 ldo_out vota ldo_in ldo_in sg13_lv_pmos L=0.5u W=8000.0u ng=1 m=1
XR2 vss pos rhigh w=0.5e-6 l=30e-6 m=1 b=0
XR1 pos ldo_out rhigh w=0.5e-6 l=10e-6 m=1 b=0
x1 vref pos iref ldo_in vss vota ota
.ends


* expanding   symbol:  xschem/ldo/ldo_openloop.sym # of pins=7
** sym_path: /home/ac3e/Documents/ihp_design/xschem/ldo/ldo_openloop.sym
** sch_path: /home/ac3e/Documents/ihp_design/xschem/ldo/ldo_openloop.sch
.subckt ldo_openloop ldo_in ldo_out iref vref vss vin_p vdiv_out
*.PININFO iref:I vin_p:I ldo_in:B vss:B vout:O vdiv_out:B ldo_out:B ldo_in:B vss:B vref:I
XM9 ldo_out vout ldo_in ldo_in sg13_lv_pmos L=0.5u W=8000.0u ng=1 m=1
XR1 vdiv_out ldo_out rhigh w=0.5e-6 l=10e-6 m=1 b=0
XR3 vss vdiv_out rhigh w=0.5e-6 l=30e-6 m=1 b=0
x1 vref vin_p iref ldo_in vss vout ota
.ends


* expanding   symbol:  xschem/pass_transistor/pass_transistor.sym # of pins=3
** sym_path: /home/ac3e/Documents/ihp_design/xschem/pass_transistor/pass_transistor.sym
** sch_path: /home/ac3e/Documents/ihp_design/xschem/pass_transistor/pass_transistor.sch
.subckt pass_transistor pt_g pt_s pt_d
*.PININFO pt_s:B pt_d:B pt_g:B
XM9 pt_d pt_g pt_s pt_s sg13_lv_pmos L=0.5u W=8000.0u ng=1 m=1
.ends


* expanding   symbol:  xschem/ota/ota.sym # of pins=6
** sym_path: /home/ac3e/Documents/ihp_design/xschem/ota/ota.sym
** sch_path: /home/ac3e/Documents/ihp_design/xschem/ota/ota.sch
.subckt ota vin_n vin_p iref vdd vss vout
*.PININFO iref:I vin_n:I vin_p:I vdd:B vss:B vout:O
XM1 net1 vin_n net2 vss sg13_lv_nmos L=2u W=15u ng=1 m=1
XM2 net3 vin_p net2 vss sg13_lv_nmos L=2u W=15u ng=1 m=1
XM3 net3 net1 vdd vdd sg13_lv_pmos L=1u W=2u ng=1 m=1
XM4 net1 net1 vdd vdd sg13_lv_pmos L=1u W=2u ng=1 m=1
XM5 net2 iref vss vss sg13_lv_nmos L=2u W=6u ng=1 m=1
XM8 iref iref vss vss sg13_lv_nmos L=2u W=6u ng=1 m=1
XM6 vout net3 vdd vdd sg13_lv_pmos L=0.5u W=20u ng=1 m=1
XM7 vout iref vss vss sg13_lv_nmos L=2u W=24u ng=1 m=1
XR2 net3 net4 rhigh w=0.5e-6 l=10e-6 m=1 b=0
XC2 vout net4 cap_cmim W=45.0e-6 L=45.0e-6 MF=1
.ends

.end